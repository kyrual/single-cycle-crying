`timescale 1ps/1ps

module mux4(A, B, C, D, Szero, Sone, Zout);
    input A, B, C, D, Szero, Sone;
    output Zout;

    wire An
endmodule